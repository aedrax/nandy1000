// Testbench
// Test   | sel  |        a         |        b         |        c         |        d         |       out        |
// Test 0 |  00  | 0000000000000000 | 0000000000000000 | 0000000000000000 | 0000000000000000 | 0000000000000000 |
// Test 1 |  01  | 0000000000000000 | 0000000000000000 | 0000000000000000 | 0000000000000000 | 0000000000000000 |
// Test 2 |  10  | 0000000000000000 | 0000000000000000 | 0000000000000000 | 0000000000000000 | 0000000000000000 |
// Test 3 |  11  | 0000000000000000 | 0000000000000000 | 0000000000000000 | 0000000000000000 | 0000000000000000 |
// Test 4 |  00  | 0001001000110100 | 1001100001110110 | 1010101010101010 | 0101010101010101 | 0001001000110100 |
// Test 5 |  01  | 0001001000110100 | 1001100001110110 | 1010101010101010 | 0101010101010101 | 1001100001110110 |
// Test 6 |  10  | 0001001000110100 | 1001100001110110 | 1010101010101010 | 0101010101010101 | 1010101010101010 |
// Test 7 |  11  | 0001001000110100 | 1001100001110110 | 1010101010101010 | 0101010101010101 | 0101010101010101 |


`include "Mux4way16bit.v"

module Mux4way16bitTest;

  reg [1:0] sel;
  reg [15:0] a;
  reg [15:0] b;
  reg [15:0] c;
  reg [15:0] d;
  wire [15:0] out;
  reg [15:0] expected;
  reg allPassed;
  
  // Instantiate design under test
  Mux4way16bit MUX4WAY16BIT(.out(out), .select(sel), .inA(a), .inB(b), .inC(c), .inD(d));

  initial begin
    // Dump waves
    $dumpfile("dump.vcd");
    $dumpvars(1);
    allPassed = 1;    
    $display("Begin Test: MUX4WAY16BIT");

    $write("Test 0: ");
    test(2'b00, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000);

    $write("Test 1: ");
    test(2'b01, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000);

    $write("Test 2: ");
    test(2'b10, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000);

    $write("Test 3: ");
    test(2'b11, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000, 16'b0000000000000000);

    $write("Test 4: ");
    test(2'b00, 16'b0001001000110100, 16'b1001100001110110, 16'b1010101010101010, 16'b0101010101010101, 16'b0001001000110100);

    $write("Test 5: ");
    test(2'b01, 16'b0001001000110100, 16'b1001100001110110, 16'b1010101010101010, 16'b0101010101010101, 16'b1001100001110110);

    $write("Test 6: ");
    test(2'b10, 16'b0001001000110100, 16'b1001100001110110, 16'b1010101010101010, 16'b0101010101010101, 16'b1010101010101010);

    $write("Test 7: ");
    test(2'b11, 16'b0001001000110100, 16'b1001100001110110, 16'b1010101010101010, 16'b0101010101010101, 16'b0101010101010101);

    
    #100
    $display("Finished Test: MUX4WAY16BIT");
    if (allPassed)
      $display("All tests PASSED");
    else
      $display("Some test has FAILED");
  end
  
  task test(input [1:0] t_sel, input [15:0] t_a, t_b, t_c, t_d, t_expected);
    sel = t_sel;
    a = t_a;
    b = t_b;
    c = t_c;
    d = t_d;
    expected = t_expected;
    #1 $write("Select:%0h, A:%0h, B:%0h, C:%0h, D:%0h, Output:%0h, Expected:%0h ", sel, a, b, c, d, out, expected);
    if (out === expected)
      $display("[PASSED]");
    else begin
      $display("[FAILED]");
      allPassed <= 0;
    end
  endtask

endmodule
